module alien(

);