module alien_laser(

);