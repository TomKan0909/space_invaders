module alien_laser(

);

// make it shoot once every 2 seconds ???