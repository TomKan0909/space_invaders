module player_laser(
    input clk,
    input reset_n,
    input shoot, // signal to shoot the laser
    input 
);